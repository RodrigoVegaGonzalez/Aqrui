module addsum();

endmodule 